
/*
 * Simple hello world example.
 * Iesus Hominum Salvator.
 */

module main;

initial
    begin
        $display("Hello, World!");
        $finish;
    end

endmodule


