
/**
 * Iesus Hominum Salvator.
 */

module supply ( output vdd, gnd );

    supply1 _vdd;
    supply0 _gnd;

    assign vdd = _vdd;
    assign gnd = _gnd;

endmodule


